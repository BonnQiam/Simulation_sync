interface intf(input logic clk,reset);
  
  //declaring the signals
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] sum;
endinterface